module and_device (a, b, s);
	input  a;
	input  b;
	output s;

	assign s = a & b;
endmodule